	component tb is
		port (
		);
	end component tb;

	u0 : component tb
		port map (
		);

