module tb (
	);
endmodule

